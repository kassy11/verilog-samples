module bgate(A, B, C, X);
  input A, B, C;
  output X;
  assign X = (A | B) & ~C;
endmodule