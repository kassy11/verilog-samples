module mux5to1(data, sw, led);
  input [4:0] data;
  output []

endmodule

module mux5to1_test();

endmodule